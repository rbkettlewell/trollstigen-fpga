
module RowDecoder ( io_rAddr, io_bAddr, io_gRows_18, io_gRows_17, io_gRows_16, 
        io_gRows_15, io_gRows_14, io_gRows_13, io_gRows_12, io_gRows_11, 
        io_gRows_10, io_gRows_9, io_gRows_8, io_gRows_7, io_gRows_6, 
        io_gRows_5, io_gRows_4, io_gRows_3, io_gRows_2, io_gRows_1, io_gRows_0
 );
  input [5:0] io_rAddr;
  input [3:0] io_bAddr;
  output [8:0] io_gRows_18;
  output [8:0] io_gRows_17;
  output [8:0] io_gRows_16;
  output [8:0] io_gRows_15;
  output [8:0] io_gRows_14;
  output [8:0] io_gRows_13;
  output [8:0] io_gRows_12;
  output [8:0] io_gRows_11;
  output [8:0] io_gRows_10;
  output [8:0] io_gRows_9;
  output [8:0] io_gRows_8;
  output [8:0] io_gRows_7;
  output [8:0] io_gRows_6;
  output [8:0] io_gRows_5;
  output [8:0] io_gRows_4;
  output [8:0] io_gRows_3;
  output [8:0] io_gRows_2;
  output [8:0] io_gRows_1;
  output [8:0] io_gRows_0;
  wire   n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504;

  INVX2TS U503 ( .A(n331), .Y(n347) );
  INVX2TS U504 ( .A(n332), .Y(n365) );
  INVX2TS U505 ( .A(n336), .Y(n337) );
  INVX2TS U506 ( .A(n333), .Y(n343) );
  INVX2TS U507 ( .A(n341), .Y(n342) );
  CLKBUFX2TS U508 ( .A(io_bAddr[1]), .Y(n330) );
  CLKBUFX2TS U509 ( .A(io_bAddr[0]), .Y(n331) );
  NOR2XLTS U510 ( .A(n330), .B(n331), .Y(n354) );
  CLKBUFX2TS U511 ( .A(n354), .Y(n398) );
  INVX2TS U512 ( .A(n398), .Y(n467) );
  CLKBUFX2TS U513 ( .A(io_rAddr[2]), .Y(n332) );
  INVX2TS U514 ( .A(n365), .Y(n413) );
  CLKBUFX2TS U515 ( .A(io_rAddr[1]), .Y(n333) );
  INVX2TS U516 ( .A(n343), .Y(n366) );
  CLKBUFX2TS U517 ( .A(io_rAddr[3]), .Y(n334) );
  INVX2TS U518 ( .A(n334), .Y(n431) );
  NAND3XLTS U519 ( .A(n365), .B(n343), .C(n431), .Y(n480) );
  CLKBUFX2TS U520 ( .A(io_rAddr[5]), .Y(n335) );
  CLKBUFX2TS U521 ( .A(io_rAddr[0]), .Y(n336) );
  CLKBUFX2TS U522 ( .A(io_rAddr[4]), .Y(n338) );
  NOR3XLTS U523 ( .A(n335), .B(n336), .C(n338), .Y(n432) );
  NAND2BXLTS U524 ( .AN(n480), .B(n432), .Y(n339) );
  INVX2TS U525 ( .A(n339), .Y(n494) );
  INVX2TS U526 ( .A(n494), .Y(n499) );
  CLKBUFX2TS U527 ( .A(io_bAddr[3]), .Y(n340) );
  CLKBUFX2TS U528 ( .A(io_bAddr[2]), .Y(n341) );
  OR2X1TS U529 ( .A(n340), .B(n341), .Y(n389) );
  INVX2TS U530 ( .A(n389), .Y(n410) );
  INVX2TS U531 ( .A(n410), .Y(n437) );
  INVX2TS U532 ( .A(n437), .Y(n395) );
  NAND2BXLTS U533 ( .AN(n499), .B(n395), .Y(n503) );
  NOR2XLTS U534 ( .A(n467), .B(n503), .Y(io_gRows_0[0]) );
  CLKAND2X2TS U535 ( .A(n366), .B(n365), .Y(n386) );
  INVX2TS U536 ( .A(n386), .Y(n456) );
  NAND3BXLTS U537 ( .AN(n335), .B(n338), .C(n337), .Y(n360) );
  NOR3XLTS U538 ( .A(n334), .B(n456), .C(n360), .Y(n351) );
  INVX2TS U539 ( .A(n351), .Y(n344) );
  CLKAND2X2TS U540 ( .A(n330), .B(n331), .Y(n370) );
  INVX2TS U541 ( .A(n370), .Y(n422) );
  INVX2TS U542 ( .A(n422), .Y(n436) );
  INVX2TS U543 ( .A(n436), .Y(n396) );
  NOR2XLTS U544 ( .A(n342), .B(n340), .Y(n349) );
  NAND2BXLTS U545 ( .AN(n396), .B(n349), .Y(n345) );
  INVX2TS U546 ( .A(n345), .Y(n402) );
  INVX2TS U547 ( .A(n402), .Y(n496) );
  NOR2XLTS U548 ( .A(n408), .B(n496), .Y(io_gRows_18[7]) );
  CLKAND2X2TS U549 ( .A(n330), .B(n347), .Y(n371) );
  INVX2TS U550 ( .A(n371), .Y(n423) );
  INVX2TS U551 ( .A(n423), .Y(n439) );
  INVX2TS U552 ( .A(n439), .Y(n397) );
  NAND2BXLTS U553 ( .AN(n397), .B(n349), .Y(n346) );
  INVX2TS U554 ( .A(n346), .Y(n403) );
  INVX2TS U555 ( .A(n403), .Y(n497) );
  NOR2XLTS U556 ( .A(n344), .B(n497), .Y(io_gRows_18[6]) );
  NOR2XLTS U557 ( .A(n347), .B(n330), .Y(n352) );
  NAND2X1TS U558 ( .A(n352), .B(n349), .Y(n348) );
  INVX2TS U559 ( .A(n348), .Y(n404) );
  INVX2TS U560 ( .A(n404), .Y(n498) );
  NOR2XLTS U561 ( .A(n408), .B(n498), .Y(io_gRows_18[5]) );
  INVX2TS U562 ( .A(n351), .Y(n408) );
  NAND2X1TS U563 ( .A(n354), .B(n349), .Y(n350) );
  INVX2TS U564 ( .A(n350), .Y(n405) );
  INVX2TS U565 ( .A(n405), .Y(n500) );
  NOR2XLTS U566 ( .A(n408), .B(n500), .Y(io_gRows_18[4]) );
  INVX2TS U567 ( .A(n370), .Y(n490) );
  INVX2TS U568 ( .A(n389), .Y(n488) );
  NAND2X1TS U569 ( .A(n488), .B(n351), .Y(n353) );
  NOR2XLTS U570 ( .A(n490), .B(n353), .Y(io_gRows_18[3]) );
  INVX2TS U571 ( .A(n371), .Y(n491) );
  NOR2XLTS U572 ( .A(n491), .B(n353), .Y(io_gRows_18[2]) );
  CLKBUFX2TS U573 ( .A(n352), .Y(n424) );
  INVX2TS U574 ( .A(n424), .Y(n492) );
  NOR2XLTS U575 ( .A(n492), .B(n353), .Y(io_gRows_18[1]) );
  INVX2TS U576 ( .A(n398), .Y(n478) );
  NOR2XLTS U577 ( .A(n478), .B(n353), .Y(io_gRows_18[0]) );
  NOR4BXLTS U578 ( .AN(n338), .B(n335), .C(n337), .D(n480), .Y(n358) );
  INVX1TS U579 ( .A(n358), .Y(n356) );
  NAND3XLTS U580 ( .A(n340), .B(n354), .C(n342), .Y(n355) );
  INVX2TS U581 ( .A(n355), .Y(n407) );
  INVX2TS U582 ( .A(n407), .Y(n495) );
  NOR2XLTS U583 ( .A(n356), .B(n495), .Y(io_gRows_17[8]) );
  INVX2TS U584 ( .A(n358), .Y(n357) );
  INVX2TS U585 ( .A(n402), .Y(n459) );
  NOR2XLTS U586 ( .A(n357), .B(n459), .Y(io_gRows_17[7]) );
  INVX2TS U587 ( .A(n403), .Y(n460) );
  NOR2XLTS U588 ( .A(n357), .B(n460), .Y(io_gRows_17[6]) );
  INVX2TS U589 ( .A(n404), .Y(n461) );
  NOR2XLTS U590 ( .A(n357), .B(n461), .Y(io_gRows_17[5]) );
  INVX2TS U591 ( .A(n405), .Y(n462) );
  NOR2XLTS U592 ( .A(n357), .B(n462), .Y(io_gRows_17[4]) );
  INVX2TS U593 ( .A(n370), .Y(n501) );
  NAND2X1TS U594 ( .A(n473), .B(n358), .Y(n359) );
  NOR2XLTS U595 ( .A(n501), .B(n359), .Y(io_gRows_17[3]) );
  INVX2TS U596 ( .A(n371), .Y(n502) );
  NOR2XLTS U597 ( .A(n502), .B(n359), .Y(io_gRows_17[2]) );
  INVX2TS U598 ( .A(n424), .Y(n504) );
  NOR2XLTS U599 ( .A(n504), .B(n359), .Y(io_gRows_17[1]) );
  INVX2TS U600 ( .A(n398), .Y(n426) );
  INVX2TS U601 ( .A(n354), .Y(n381) );
  NOR2XLTS U602 ( .A(n381), .B(n359), .Y(io_gRows_17[0]) );
  NOR2XLTS U603 ( .A(n360), .B(n480), .Y(n363) );
  INVX2TS U604 ( .A(n363), .Y(n361) );
  INVX2TS U605 ( .A(n407), .Y(n458) );
  NOR2XLTS U606 ( .A(n361), .B(n458), .Y(io_gRows_16[8]) );
  INVX2TS U607 ( .A(n363), .Y(n362) );
  NOR2XLTS U608 ( .A(n362), .B(n459), .Y(io_gRows_16[7]) );
  NOR2XLTS U609 ( .A(n362), .B(n460), .Y(io_gRows_16[6]) );
  NOR2XLTS U610 ( .A(n362), .B(n461), .Y(io_gRows_16[5]) );
  NOR2XLTS U611 ( .A(n362), .B(n462), .Y(io_gRows_16[4]) );
  NAND2X1TS U612 ( .A(n395), .B(n363), .Y(n364) );
  NOR2XLTS U613 ( .A(n422), .B(n364), .Y(io_gRows_16[3]) );
  NOR2XLTS U614 ( .A(n423), .B(n364), .Y(io_gRows_16[2]) );
  INVX2TS U615 ( .A(n424), .Y(n440) );
  NOR2XLTS U616 ( .A(n465), .B(n364), .Y(io_gRows_16[1]) );
  NOR2XLTS U617 ( .A(n467), .B(n364), .Y(io_gRows_16[0]) );
  NAND2X1TS U618 ( .A(n413), .B(n366), .Y(n433) );
  NOR3XLTS U619 ( .A(n335), .B(n338), .C(n337), .Y(n479) );
  NAND2X1TS U620 ( .A(n334), .B(n479), .Y(n400) );
  NOR2XLTS U621 ( .A(n433), .B(n400), .Y(n369) );
  INVX2TS U622 ( .A(n369), .Y(n367) );
  NOR2XLTS U623 ( .A(n367), .B(n458), .Y(io_gRows_15[8]) );
  INVX2TS U624 ( .A(n369), .Y(n368) );
  INVX2TS U625 ( .A(n402), .Y(n416) );
  NOR2XLTS U626 ( .A(n368), .B(n416), .Y(io_gRows_15[7]) );
  INVX2TS U627 ( .A(n403), .Y(n417) );
  NOR2XLTS U628 ( .A(n368), .B(n417), .Y(io_gRows_15[6]) );
  INVX2TS U629 ( .A(n404), .Y(n418) );
  NOR2XLTS U630 ( .A(n368), .B(n418), .Y(io_gRows_15[5]) );
  INVX2TS U631 ( .A(n405), .Y(n419) );
  NOR2XLTS U632 ( .A(n368), .B(n419), .Y(io_gRows_15[4]) );
  NAND2X1TS U633 ( .A(n410), .B(n369), .Y(n372) );
  INVX2TS U634 ( .A(n370), .Y(n451) );
  NOR2XLTS U635 ( .A(n372), .B(n451), .Y(io_gRows_15[3]) );
  INVX2TS U636 ( .A(n371), .Y(n452) );
  NOR2XLTS U637 ( .A(n372), .B(n452), .Y(io_gRows_15[2]) );
  NOR2XLTS U638 ( .A(n372), .B(n476), .Y(io_gRows_15[1]) );
  NOR2XLTS U639 ( .A(n478), .B(n372), .Y(io_gRows_15[0]) );
  NAND2X1TS U640 ( .A(n334), .B(n432), .Y(n412) );
  NOR2XLTS U641 ( .A(n433), .B(n412), .Y(n375) );
  INVX2TS U642 ( .A(n375), .Y(n373) );
  INVX2TS U643 ( .A(n407), .Y(n414) );
  NOR2XLTS U644 ( .A(n373), .B(n414), .Y(io_gRows_14[8]) );
  INVX2TS U645 ( .A(n375), .Y(n374) );
  NOR2XLTS U646 ( .A(n374), .B(n496), .Y(io_gRows_14[7]) );
  NOR2XLTS U647 ( .A(n374), .B(n497), .Y(io_gRows_14[6]) );
  NOR2XLTS U648 ( .A(n374), .B(n498), .Y(io_gRows_14[5]) );
  NOR2XLTS U649 ( .A(n374), .B(n500), .Y(io_gRows_14[4]) );
  NAND2X1TS U650 ( .A(n395), .B(n375), .Y(n376) );
  NOR2XLTS U651 ( .A(n396), .B(n376), .Y(io_gRows_14[3]) );
  NOR2XLTS U652 ( .A(n397), .B(n376), .Y(io_gRows_14[2]) );
  NOR2XLTS U653 ( .A(n492), .B(n376), .Y(io_gRows_14[1]) );
  NOR2XLTS U654 ( .A(n426), .B(n376), .Y(io_gRows_14[0]) );
  NAND2X1TS U655 ( .A(n332), .B(n343), .Y(n447) );
  NOR2XLTS U656 ( .A(n400), .B(n447), .Y(n379) );
  INVX2TS U657 ( .A(n379), .Y(n377) );
  NOR2XLTS U658 ( .A(n377), .B(n495), .Y(io_gRows_13[8]) );
  INVX2TS U659 ( .A(n379), .Y(n378) );
  NOR2XLTS U660 ( .A(n378), .B(n345), .Y(io_gRows_13[7]) );
  NOR2XLTS U661 ( .A(n378), .B(n346), .Y(io_gRows_13[6]) );
  NOR2XLTS U662 ( .A(n378), .B(n348), .Y(io_gRows_13[5]) );
  NOR2XLTS U663 ( .A(n378), .B(n350), .Y(io_gRows_13[4]) );
  NAND2X1TS U664 ( .A(n445), .B(n379), .Y(n380) );
  NOR2XLTS U665 ( .A(n422), .B(n380), .Y(io_gRows_13[3]) );
  NOR2XLTS U666 ( .A(n423), .B(n380), .Y(io_gRows_13[2]) );
  NOR2XLTS U667 ( .A(n504), .B(n380), .Y(io_gRows_13[1]) );
  NOR2XLTS U668 ( .A(n381), .B(n380), .Y(io_gRows_13[0]) );
  NOR2XLTS U669 ( .A(n412), .B(n447), .Y(n384) );
  INVX2TS U670 ( .A(n384), .Y(n382) );
  NOR2XLTS U671 ( .A(n382), .B(n355), .Y(io_gRows_12[8]) );
  INVX2TS U672 ( .A(n384), .Y(n383) );
  NOR2XLTS U673 ( .A(n383), .B(n416), .Y(io_gRows_12[7]) );
  NOR2XLTS U674 ( .A(n383), .B(n417), .Y(io_gRows_12[6]) );
  NOR2XLTS U675 ( .A(n383), .B(n418), .Y(io_gRows_12[5]) );
  NOR2XLTS U676 ( .A(n383), .B(n419), .Y(io_gRows_12[4]) );
  NAND2X1TS U677 ( .A(n410), .B(n384), .Y(n385) );
  NOR2XLTS U678 ( .A(n490), .B(n385), .Y(io_gRows_12[3]) );
  NOR2XLTS U679 ( .A(n491), .B(n385), .Y(io_gRows_12[2]) );
  NOR2XLTS U680 ( .A(n440), .B(n385), .Y(io_gRows_12[1]) );
  NOR2XLTS U681 ( .A(n478), .B(n385), .Y(io_gRows_12[0]) );
  INVX2TS U682 ( .A(n386), .Y(n469) );
  NOR2XLTS U683 ( .A(n400), .B(n469), .Y(n390) );
  INVX2TS U684 ( .A(n390), .Y(n387) );
  NOR2XLTS U685 ( .A(n388), .B(n414), .Y(io_gRows_11[8]) );
  NOR2XLTS U686 ( .A(n387), .B(n459), .Y(io_gRows_11[7]) );
  NOR2XLTS U687 ( .A(n388), .B(n460), .Y(io_gRows_11[6]) );
  INVX2TS U688 ( .A(n390), .Y(n388) );
  NOR2XLTS U689 ( .A(n388), .B(n461), .Y(io_gRows_11[5]) );
  NOR2XLTS U690 ( .A(n388), .B(n462), .Y(io_gRows_11[4]) );
  INVX2TS U691 ( .A(n389), .Y(n445) );
  NAND2X1TS U692 ( .A(n445), .B(n390), .Y(n391) );
  NOR2XLTS U693 ( .A(n451), .B(n391), .Y(io_gRows_11[3]) );
  NOR2XLTS U694 ( .A(n452), .B(n391), .Y(io_gRows_11[2]) );
  NOR2XLTS U695 ( .A(n465), .B(n391), .Y(io_gRows_11[1]) );
  NOR2XLTS U696 ( .A(n426), .B(n391), .Y(io_gRows_11[0]) );
  NOR2XLTS U697 ( .A(n412), .B(n456), .Y(n394) );
  INVX2TS U698 ( .A(n394), .Y(n392) );
  NOR2XLTS U699 ( .A(n393), .B(n458), .Y(io_gRows_10[8]) );
  NOR2XLTS U700 ( .A(n392), .B(n345), .Y(io_gRows_10[7]) );
  NOR2XLTS U701 ( .A(n393), .B(n346), .Y(io_gRows_10[6]) );
  INVX2TS U702 ( .A(n394), .Y(n393) );
  NOR2XLTS U703 ( .A(n393), .B(n348), .Y(io_gRows_10[5]) );
  NOR2XLTS U704 ( .A(n393), .B(n350), .Y(io_gRows_10[4]) );
  NAND2X1TS U705 ( .A(n395), .B(n394), .Y(n399) );
  NOR2XLTS U706 ( .A(n396), .B(n399), .Y(io_gRows_10[3]) );
  NOR2XLTS U707 ( .A(n397), .B(n399), .Y(io_gRows_10[2]) );
  NOR2XLTS U708 ( .A(n504), .B(n399), .Y(io_gRows_10[1]) );
  INVX2TS U709 ( .A(n398), .Y(n454) );
  NOR2XLTS U710 ( .A(n454), .B(n399), .Y(io_gRows_10[0]) );
  NOR3XLTS U711 ( .A(n413), .B(n333), .C(n400), .Y(n409) );
  INVX2TS U712 ( .A(n409), .Y(n401) );
  NOR2XLTS U713 ( .A(n401), .B(n355), .Y(io_gRows_9[8]) );
  INVX2TS U714 ( .A(n409), .Y(n406) );
  INVX2TS U715 ( .A(n402), .Y(n483) );
  NOR2XLTS U716 ( .A(n406), .B(n483), .Y(io_gRows_9[7]) );
  INVX2TS U717 ( .A(n403), .Y(n484) );
  NOR2XLTS U718 ( .A(n406), .B(n484), .Y(io_gRows_9[6]) );
  INVX2TS U719 ( .A(n404), .Y(n486) );
  NOR2XLTS U720 ( .A(n406), .B(n486), .Y(io_gRows_9[5]) );
  INVX2TS U721 ( .A(n405), .Y(n487) );
  NOR2XLTS U722 ( .A(n406), .B(n487), .Y(io_gRows_9[4]) );
  INVX2TS U723 ( .A(n407), .Y(n482) );
  NOR2XLTS U724 ( .A(n408), .B(n482), .Y(io_gRows_18[8]) );
  NAND2X1TS U725 ( .A(n410), .B(n409), .Y(n411) );
  NOR2XLTS U726 ( .A(n451), .B(n411), .Y(io_gRows_9[3]) );
  NOR2XLTS U727 ( .A(n452), .B(n411), .Y(io_gRows_9[2]) );
  NOR2XLTS U728 ( .A(n440), .B(n411), .Y(io_gRows_9[1]) );
  NOR2XLTS U729 ( .A(n381), .B(n411), .Y(io_gRows_9[0]) );
  NOR3XLTS U730 ( .A(n413), .B(n366), .C(n412), .Y(n421) );
  INVX2TS U731 ( .A(n421), .Y(n415) );
  NOR2XLTS U732 ( .A(n415), .B(n414), .Y(io_gRows_8[8]) );
  INVX2TS U733 ( .A(n421), .Y(n420) );
  NOR2XLTS U734 ( .A(n420), .B(n416), .Y(io_gRows_8[7]) );
  NOR2XLTS U735 ( .A(n420), .B(n417), .Y(io_gRows_8[6]) );
  NOR2XLTS U736 ( .A(n420), .B(n418), .Y(io_gRows_8[5]) );
  NOR2XLTS U737 ( .A(n420), .B(n419), .Y(io_gRows_8[4]) );
  NAND2X1TS U738 ( .A(n445), .B(n421), .Y(n425) );
  NOR2XLTS U739 ( .A(n422), .B(n425), .Y(io_gRows_8[3]) );
  NOR2XLTS U740 ( .A(n423), .B(n425), .Y(io_gRows_8[2]) );
  INVX2TS U741 ( .A(n424), .Y(n476) );
  NOR2XLTS U742 ( .A(n476), .B(n425), .Y(io_gRows_8[1]) );
  NOR2XLTS U743 ( .A(n426), .B(n425), .Y(io_gRows_8[0]) );
  NAND2X1TS U744 ( .A(n479), .B(n431), .Y(n455) );
  NOR2XLTS U745 ( .A(n433), .B(n455), .Y(n429) );
  INVX2TS U746 ( .A(n429), .Y(n427) );
  NOR2XLTS U747 ( .A(n427), .B(n355), .Y(io_gRows_7[8]) );
  INVX2TS U748 ( .A(n429), .Y(n428) );
  NOR2XLTS U749 ( .A(n428), .B(n345), .Y(io_gRows_7[7]) );
  NOR2XLTS U750 ( .A(n428), .B(n346), .Y(io_gRows_7[6]) );
  NOR2XLTS U751 ( .A(n428), .B(n348), .Y(io_gRows_7[5]) );
  NOR2XLTS U752 ( .A(n428), .B(n350), .Y(io_gRows_7[4]) );
  NAND2X1TS U753 ( .A(n488), .B(n429), .Y(n430) );
  NOR2XLTS U754 ( .A(n501), .B(n430), .Y(io_gRows_7[3]) );
  NOR2XLTS U755 ( .A(n502), .B(n430), .Y(io_gRows_7[2]) );
  INVX2TS U756 ( .A(n352), .Y(n465) );
  NOR2XLTS U757 ( .A(n465), .B(n430), .Y(io_gRows_7[1]) );
  NOR2XLTS U758 ( .A(n454), .B(n430), .Y(io_gRows_7[0]) );
  NAND2X1TS U759 ( .A(n432), .B(n431), .Y(n468) );
  NOR2XLTS U760 ( .A(n433), .B(n468), .Y(n438) );
  INVX2TS U761 ( .A(n438), .Y(n434) );
  NOR2XLTS U762 ( .A(n434), .B(n495), .Y(io_gRows_6[8]) );
  INVX2TS U763 ( .A(n438), .Y(n435) );
  NOR2XLTS U764 ( .A(n435), .B(n496), .Y(io_gRows_6[7]) );
  NOR2XLTS U765 ( .A(n435), .B(n497), .Y(io_gRows_6[6]) );
  NOR2XLTS U766 ( .A(n435), .B(n498), .Y(io_gRows_6[5]) );
  NOR2XLTS U767 ( .A(n435), .B(n500), .Y(io_gRows_6[4]) );
  INVX2TS U768 ( .A(n436), .Y(n474) );
  INVX2TS U769 ( .A(n437), .Y(n473) );
  NAND2X1TS U770 ( .A(n473), .B(n438), .Y(n441) );
  NOR2XLTS U771 ( .A(n474), .B(n441), .Y(io_gRows_6[3]) );
  INVX2TS U772 ( .A(n439), .Y(n475) );
  NOR2XLTS U773 ( .A(n475), .B(n441), .Y(io_gRows_6[2]) );
  NOR2XLTS U774 ( .A(n440), .B(n441), .Y(io_gRows_6[1]) );
  NOR2XLTS U775 ( .A(n467), .B(n441), .Y(io_gRows_6[0]) );
  NOR2XLTS U776 ( .A(n447), .B(n455), .Y(n444) );
  INVX2TS U777 ( .A(n444), .Y(n442) );
  NOR2XLTS U778 ( .A(n442), .B(n482), .Y(io_gRows_5[8]) );
  INVX2TS U779 ( .A(n444), .Y(n443) );
  NOR2XLTS U780 ( .A(n443), .B(n483), .Y(io_gRows_5[7]) );
  NOR2XLTS U781 ( .A(n443), .B(n484), .Y(io_gRows_5[6]) );
  NOR2XLTS U782 ( .A(n443), .B(n486), .Y(io_gRows_5[5]) );
  NOR2XLTS U783 ( .A(n443), .B(n487), .Y(io_gRows_5[4]) );
  NAND2X1TS U784 ( .A(n445), .B(n444), .Y(n446) );
  NOR2XLTS U785 ( .A(n501), .B(n446), .Y(io_gRows_5[3]) );
  NOR2XLTS U786 ( .A(n502), .B(n446), .Y(io_gRows_5[2]) );
  NOR2XLTS U787 ( .A(n476), .B(n446), .Y(io_gRows_5[1]) );
  NOR2XLTS U788 ( .A(n381), .B(n446), .Y(io_gRows_5[0]) );
  NOR2XLTS U789 ( .A(n447), .B(n468), .Y(n450) );
  INVX2TS U790 ( .A(n450), .Y(n448) );
  NOR2XLTS U791 ( .A(n448), .B(n414), .Y(io_gRows_4[8]) );
  INVX2TS U792 ( .A(n450), .Y(n449) );
  NOR2XLTS U793 ( .A(n449), .B(n416), .Y(io_gRows_4[7]) );
  NOR2XLTS U794 ( .A(n449), .B(n417), .Y(io_gRows_4[6]) );
  NOR2XLTS U795 ( .A(n449), .B(n418), .Y(io_gRows_4[5]) );
  NOR2XLTS U796 ( .A(n449), .B(n419), .Y(io_gRows_4[4]) );
  NAND2X1TS U797 ( .A(n488), .B(n450), .Y(n453) );
  NOR2XLTS U798 ( .A(n451), .B(n453), .Y(io_gRows_4[3]) );
  NOR2XLTS U799 ( .A(n452), .B(n453), .Y(io_gRows_4[2]) );
  NOR2XLTS U800 ( .A(n492), .B(n453), .Y(io_gRows_4[1]) );
  NOR2XLTS U801 ( .A(n454), .B(n453), .Y(io_gRows_4[0]) );
  NOR2XLTS U802 ( .A(n456), .B(n455), .Y(n464) );
  INVX2TS U803 ( .A(n464), .Y(n457) );
  NOR2XLTS U804 ( .A(n463), .B(n458), .Y(io_gRows_3[8]) );
  NOR2XLTS U805 ( .A(n457), .B(n459), .Y(io_gRows_3[7]) );
  NOR2XLTS U806 ( .A(n463), .B(n460), .Y(io_gRows_3[6]) );
  INVX2TS U807 ( .A(n464), .Y(n463) );
  NOR2XLTS U808 ( .A(n463), .B(n461), .Y(io_gRows_3[5]) );
  NOR2XLTS U809 ( .A(n463), .B(n462), .Y(io_gRows_3[4]) );
  NAND2X1TS U810 ( .A(n473), .B(n464), .Y(n466) );
  NOR2XLTS U811 ( .A(n490), .B(n466), .Y(io_gRows_3[3]) );
  NOR2XLTS U812 ( .A(n491), .B(n466), .Y(io_gRows_3[2]) );
  NOR2XLTS U813 ( .A(n465), .B(n466), .Y(io_gRows_3[1]) );
  NOR2XLTS U814 ( .A(n467), .B(n466), .Y(io_gRows_3[0]) );
  NOR2XLTS U815 ( .A(n469), .B(n468), .Y(n472) );
  INVX2TS U816 ( .A(n472), .Y(n470) );
  NOR2XLTS U817 ( .A(n471), .B(n482), .Y(io_gRows_2[8]) );
  NOR2XLTS U818 ( .A(n470), .B(n483), .Y(io_gRows_2[7]) );
  NOR2XLTS U819 ( .A(n471), .B(n484), .Y(io_gRows_2[6]) );
  INVX2TS U820 ( .A(n472), .Y(n471) );
  NOR2XLTS U821 ( .A(n471), .B(n486), .Y(io_gRows_2[5]) );
  NOR2XLTS U822 ( .A(n471), .B(n487), .Y(io_gRows_2[4]) );
  NAND2X1TS U823 ( .A(n473), .B(n472), .Y(n477) );
  NOR2XLTS U824 ( .A(n474), .B(n477), .Y(io_gRows_2[3]) );
  NOR2XLTS U825 ( .A(n475), .B(n477), .Y(io_gRows_2[2]) );
  NOR2XLTS U826 ( .A(n476), .B(n477), .Y(io_gRows_2[1]) );
  NOR2XLTS U827 ( .A(n478), .B(n477), .Y(io_gRows_2[0]) );
  NAND2BXLTS U828 ( .AN(n480), .B(n479), .Y(n481) );
  INVX2TS U829 ( .A(n481), .Y(n485) );
  NOR2XLTS U830 ( .A(n482), .B(n481), .Y(io_gRows_1[8]) );
  NOR2XLTS U831 ( .A(n483), .B(n489), .Y(io_gRows_1[7]) );
  NOR2XLTS U832 ( .A(n484), .B(n481), .Y(io_gRows_1[6]) );
  INVX2TS U833 ( .A(n485), .Y(n489) );
  NOR2XLTS U834 ( .A(n486), .B(n489), .Y(io_gRows_1[5]) );
  NOR2XLTS U835 ( .A(n487), .B(n489), .Y(io_gRows_1[4]) );
  NAND2BXLTS U836 ( .AN(n489), .B(n488), .Y(n493) );
  NOR2XLTS U837 ( .A(n490), .B(n493), .Y(io_gRows_1[3]) );
  NOR2XLTS U838 ( .A(n491), .B(n493), .Y(io_gRows_1[2]) );
  NOR2XLTS U839 ( .A(n492), .B(n493), .Y(io_gRows_1[1]) );
  NOR2XLTS U840 ( .A(n454), .B(n493), .Y(io_gRows_1[0]) );
  NOR2XLTS U841 ( .A(n495), .B(n339), .Y(io_gRows_0[8]) );
  NOR2XLTS U842 ( .A(n496), .B(n499), .Y(io_gRows_0[7]) );
  NOR2XLTS U843 ( .A(n497), .B(n339), .Y(io_gRows_0[6]) );
  NOR2XLTS U844 ( .A(n498), .B(n499), .Y(io_gRows_0[5]) );
  NOR2XLTS U845 ( .A(n500), .B(n499), .Y(io_gRows_0[4]) );
  NOR2XLTS U846 ( .A(n501), .B(n503), .Y(io_gRows_0[3]) );
  NOR2XLTS U847 ( .A(n502), .B(n503), .Y(io_gRows_0[2]) );
  NOR2XLTS U848 ( .A(n504), .B(n503), .Y(io_gRows_0[1]) );
endmodule

