
module ColumnDecoder ( io_WE, io_RE, io_bRead, io_bWrite, io_byteRead_14, 
        io_byteRead_13, io_byteRead_12, io_byteRead_11, io_byteRead_10, 
        io_byteRead_9, io_byteRead_8, io_byteRead_7, io_byteRead_6, 
        io_byteRead_5, io_byteRead_4, io_byteRead_3, io_byteRead_2, 
        io_byteRead_1, io_byteRead_0, io_byteWrite_14, io_byteWrite_13, 
        io_byteWrite_12, io_byteWrite_11, io_byteWrite_10, io_byteWrite_9, 
        io_byteWrite_8, io_byteWrite_7, io_byteWrite_6, io_byteWrite_5, 
        io_byteWrite_4, io_byteWrite_3, io_byteWrite_2, io_byteWrite_1, 
        io_byteWrite_0, io_cAddr, io_cDataIn, io_cDataOut );
  output [14:0] io_bRead;
  output [14:0] io_bWrite;
  input [0:7] io_byteRead_14;
  input [0:7] io_byteRead_13;
  input [0:7] io_byteRead_12;
  input [0:7] io_byteRead_11;
  input [0:7] io_byteRead_10;
  input [0:7] io_byteRead_9;
  input [0:7] io_byteRead_8;
  input [0:7] io_byteRead_7;
  input [0:7] io_byteRead_6;
  input [0:7] io_byteRead_5;
  input [0:7] io_byteRead_4;
  input [0:7] io_byteRead_3;
  input [0:7] io_byteRead_2;
  input [0:7] io_byteRead_1;
  input [0:7] io_byteRead_0;
  output [0:7] io_byteWrite_14;
  output [0:7] io_byteWrite_13;
  output [0:7] io_byteWrite_12;
  output [0:7] io_byteWrite_11;
  output [0:7] io_byteWrite_10;
  output [0:7] io_byteWrite_9;
  output [0:7] io_byteWrite_8;
  output [0:7] io_byteWrite_7;
  output [0:7] io_byteWrite_6;
  output [0:7] io_byteWrite_5;
  output [0:7] io_byteWrite_4;
  output [0:7] io_byteWrite_3;
  output [0:7] io_byteWrite_2;
  output [0:7] io_byteWrite_1;
  output [0:7] io_byteWrite_0;
  input [3:0] io_cAddr;
  input [7:0] io_cDataIn;
  output [7:0] io_cDataOut;
  input io_WE, io_RE;
  wire   n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n475, n477,
         n479, n481, n483, n485, n487, n489, n491, n493, n495, n496, n498,
         n500, n502, n504, n505, n506, n507, n508, n509, n510, n511, n512;
  wire   [0:7] io_cDataInBigEndian;
  assign io_cDataInBigEndian[0] = io_cDataIn[0];
  assign io_cDataInBigEndian[1] = io_cDataIn[1];
  assign io_cDataInBigEndian[2] = io_cDataIn[2];
  assign io_cDataInBigEndian[3] = io_cDataIn[3];
  assign io_cDataInBigEndian[4] = io_cDataIn[4];
  assign io_cDataInBigEndian[5] = io_cDataIn[5];
  assign io_cDataInBigEndian[6] = io_cDataIn[6];
  assign io_cDataInBigEndian[7] = io_cDataIn[7];

  TLATXLTS \io_cDataInBigEndianLatched_reg[0]  ( .G(n495), .D(
        io_cDataInBigEndian[0]), .Q(io_byteWrite_1[0]), .QN(n512) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[1]  ( .G(n496), .D(
        io_cDataInBigEndian[1]), .Q(io_byteWrite_1[1]), .QN(n511) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[2]  ( .G(n496), .D(
        io_cDataInBigEndian[2]), .Q(io_byteWrite_1[2]), .QN(n510) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[3]  ( .G(n495), .D(
        io_cDataInBigEndian[3]), .Q(io_byteWrite_1[3]), .QN(n509) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[4]  ( .G(n294), .D(
        io_cDataInBigEndian[4]), .Q(io_byteWrite_1[4]), .QN(n508) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[5]  ( .G(n496), .D(
        io_cDataInBigEndian[5]), .Q(io_byteWrite_1[5]), .QN(n507) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[6]  ( .G(n495), .D(
        io_cDataInBigEndian[6]), .Q(io_byteWrite_1[6]), .QN(n506) );
  TLATXLTS \io_cDataInBigEndianLatched_reg[7]  ( .G(n294), .D(
        io_cDataInBigEndian[7]), .Q(io_byteWrite_1[7]), .QN(n505) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[7]  ( .A(n305), .OE(n498), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[6]  ( .A(n306), .OE(io_bRead[0]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[5]  ( .A(n307), .OE(n498), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[4]  ( .A(n308), .OE(io_bRead[0]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[3]  ( .A(n309), .OE(n498), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[2]  ( .A(n310), .OE(io_bRead[0]), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[1]  ( .A(n311), .OE(n498), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri15[0]  ( .A(n312), .OE(io_bRead[0]), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[7]  ( .A(n313), .OE(io_bRead[1]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[6]  ( .A(n314), .OE(io_bRead[1]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[5]  ( .A(n315), .OE(io_bRead[1]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[4]  ( .A(n316), .OE(io_bRead[1]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[3]  ( .A(n317), .OE(n473), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[2]  ( .A(n318), .OE(n473), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[1]  ( .A(n319), .OE(n473), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri14[0]  ( .A(n320), .OE(n473), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[7]  ( .A(n321), .OE(io_bRead[2]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[6]  ( .A(n322), .OE(io_bRead[2]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[5]  ( .A(n323), .OE(io_bRead[2]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[4]  ( .A(n324), .OE(io_bRead[2]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[3]  ( .A(n325), .OE(n475), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[2]  ( .A(n326), .OE(n475), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[1]  ( .A(n327), .OE(n475), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri13[0]  ( .A(n328), .OE(n475), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[7]  ( .A(n329), .OE(n500), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[6]  ( .A(n330), .OE(io_bRead[3]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[5]  ( .A(n331), .OE(n500), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[4]  ( .A(n332), .OE(io_bRead[3]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[3]  ( .A(n333), .OE(n500), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[2]  ( .A(n334), .OE(io_bRead[3]), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[1]  ( .A(n335), .OE(n500), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri12[0]  ( .A(n336), .OE(io_bRead[3]), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[7]  ( .A(n337), .OE(io_bRead[4]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[6]  ( .A(n338), .OE(io_bRead[4]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[5]  ( .A(n339), .OE(io_bRead[4]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[4]  ( .A(n340), .OE(io_bRead[4]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[3]  ( .A(n341), .OE(n477), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[2]  ( .A(n342), .OE(n477), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[1]  ( .A(n343), .OE(n477), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri11[0]  ( .A(n344), .OE(n477), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[7]  ( .A(n345), .OE(io_bRead[5]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[6]  ( .A(n346), .OE(io_bRead[5]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[5]  ( .A(n347), .OE(io_bRead[5]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[4]  ( .A(n348), .OE(io_bRead[5]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[3]  ( .A(n349), .OE(n479), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[2]  ( .A(n350), .OE(n479), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[1]  ( .A(n351), .OE(n479), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri10[0]  ( .A(n352), .OE(n479), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[7]  ( .A(n353), .OE(io_bRead[6]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[6]  ( .A(n354), .OE(io_bRead[6]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[5]  ( .A(n355), .OE(io_bRead[6]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[4]  ( .A(n356), .OE(io_bRead[6]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[3]  ( .A(n357), .OE(n481), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[2]  ( .A(n358), .OE(n481), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[1]  ( .A(n359), .OE(n481), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri9[0]  ( .A(n360), .OE(n481), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[7]  ( .A(n361), .OE(io_bRead[7]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[6]  ( .A(n362), .OE(io_bRead[7]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[5]  ( .A(n363), .OE(io_bRead[7]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[4]  ( .A(n364), .OE(io_bRead[7]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[3]  ( .A(n365), .OE(n483), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[2]  ( .A(n366), .OE(n483), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[1]  ( .A(n367), .OE(n483), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri8[0]  ( .A(n368), .OE(n483), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[7]  ( .A(n369), .OE(io_bRead[8]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[6]  ( .A(n370), .OE(io_bRead[8]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[5]  ( .A(n371), .OE(io_bRead[8]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[4]  ( .A(n372), .OE(io_bRead[8]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[3]  ( .A(n373), .OE(n485), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[2]  ( .A(n374), .OE(n485), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[1]  ( .A(n375), .OE(n485), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri7[0]  ( .A(n376), .OE(n485), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[7]  ( .A(n377), .OE(io_bRead[9]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[6]  ( .A(n378), .OE(io_bRead[9]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[5]  ( .A(n379), .OE(io_bRead[9]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[4]  ( .A(n380), .OE(io_bRead[9]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[3]  ( .A(n381), .OE(n487), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[2]  ( .A(n382), .OE(n487), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[1]  ( .A(n383), .OE(n487), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri6[0]  ( .A(n384), .OE(n487), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[7]  ( .A(n385), .OE(io_bRead[10]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[6]  ( .A(n386), .OE(io_bRead[10]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[5]  ( .A(n387), .OE(io_bRead[10]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[4]  ( .A(n388), .OE(io_bRead[10]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[3]  ( .A(n389), .OE(n489), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[2]  ( .A(n390), .OE(n489), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[1]  ( .A(n391), .OE(n489), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri5[0]  ( .A(n392), .OE(n489), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[7]  ( .A(n393), .OE(io_bRead[11]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[6]  ( .A(n394), .OE(io_bRead[11]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[5]  ( .A(n395), .OE(io_bRead[11]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[4]  ( .A(n396), .OE(io_bRead[11]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[3]  ( .A(n397), .OE(n491), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[2]  ( .A(n398), .OE(n491), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[1]  ( .A(n399), .OE(n491), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri4[0]  ( .A(n400), .OE(n491), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[7]  ( .A(n401), .OE(io_bRead[12]), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[6]  ( .A(n402), .OE(io_bRead[12]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[5]  ( .A(n403), .OE(io_bRead[12]), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[4]  ( .A(n404), .OE(io_bRead[12]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[3]  ( .A(n405), .OE(n493), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[2]  ( .A(n406), .OE(n493), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[1]  ( .A(n407), .OE(n493), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri3[0]  ( .A(n408), .OE(n493), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[7]  ( .A(n409), .OE(n502), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[6]  ( .A(n410), .OE(io_bRead[13]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[5]  ( .A(n411), .OE(n502), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[4]  ( .A(n412), .OE(io_bRead[13]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[3]  ( .A(n413), .OE(n502), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[2]  ( .A(n414), .OE(io_bRead[13]), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[1]  ( .A(n415), .OE(n502), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri2[0]  ( .A(n416), .OE(io_bRead[13]), .Y(
        io_cDataOut[0]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[7]  ( .A(n417), .OE(n504), .Y(
        io_cDataOut[7]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[6]  ( .A(n418), .OE(io_bRead[14]), .Y(
        io_cDataOut[6]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[5]  ( .A(n419), .OE(n504), .Y(
        io_cDataOut[5]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[4]  ( .A(n420), .OE(io_bRead[14]), .Y(
        io_cDataOut[4]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[3]  ( .A(n421), .OE(n504), .Y(
        io_cDataOut[3]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[2]  ( .A(n422), .OE(io_bRead[14]), .Y(
        io_cDataOut[2]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[1]  ( .A(n423), .OE(n504), .Y(
        io_cDataOut[1]) );
  TBUFX2TS \io_cDataOutBigEndian_tri[0]  ( .A(n424), .OE(io_bRead[14]), .Y(
        io_cDataOut[0]) );
  NOR2XLTS U85 ( .A(n292), .B(n295), .Y(n437) );
  NAND2BXLTS U86 ( .AN(n290), .B(n291), .Y(n296) );
  NAND2BXLTS U87 ( .AN(n291), .B(n290), .Y(n299) );
  NAND4XLTS U88 ( .A(n302), .B(n303), .C(n293), .D(n304), .Y(n432) );
  NAND4XLTS U89 ( .A(n303), .B(n293), .C(n304), .D(n297), .Y(n435) );
  NAND4XLTS U90 ( .A(n302), .B(n293), .C(n304), .D(n298), .Y(n429) );
  NAND3XLTS U91 ( .A(n437), .B(n293), .C(n304), .Y(n426) );
  INVX2TS U92 ( .A(n449), .Y(io_byteWrite_0[7]) );
  INVX2TS U93 ( .A(n472), .Y(io_byteWrite_5[6]) );
  INVX2TS U94 ( .A(n471), .Y(io_byteWrite_5[5]) );
  INVX2TS U95 ( .A(n470), .Y(io_byteWrite_5[4]) );
  INVX2TS U96 ( .A(n469), .Y(io_byteWrite_5[3]) );
  INVX2TS U97 ( .A(n468), .Y(io_byteWrite_5[2]) );
  INVX2TS U98 ( .A(n467), .Y(io_byteWrite_5[1]) );
  INVX2TS U99 ( .A(n466), .Y(io_byteWrite_5[0]) );
  INVX2TS U100 ( .A(n465), .Y(io_byteWrite_6[7]) );
  INVX2TS U101 ( .A(n464), .Y(io_byteWrite_6[6]) );
  INVX2TS U102 ( .A(n463), .Y(io_byteWrite_6[5]) );
  INVX2TS U103 ( .A(n462), .Y(io_byteWrite_6[4]) );
  INVX2TS U104 ( .A(n461), .Y(io_byteWrite_6[3]) );
  INVX2TS U105 ( .A(n460), .Y(io_byteWrite_6[2]) );
  INVX2TS U106 ( .A(n459), .Y(io_byteWrite_6[1]) );
  INVX2TS U107 ( .A(n458), .Y(io_byteWrite_6[0]) );
  INVX2TS U108 ( .A(n457), .Y(io_byteWrite_7[7]) );
  INVX2TS U109 ( .A(n456), .Y(io_byteWrite_7[6]) );
  INVX2TS U110 ( .A(n455), .Y(io_byteWrite_7[5]) );
  INVX2TS U111 ( .A(n454), .Y(io_byteWrite_7[4]) );
  INVX2TS U112 ( .A(n453), .Y(io_byteWrite_7[3]) );
  INVX2TS U113 ( .A(n452), .Y(io_byteWrite_7[2]) );
  INVX2TS U114 ( .A(n451), .Y(io_byteWrite_7[1]) );
  INVX2TS U115 ( .A(n450), .Y(io_byteWrite_7[0]) );
  INVX2TS U116 ( .A(n449), .Y(io_byteWrite_8[7]) );
  INVX2TS U117 ( .A(n472), .Y(io_byteWrite_8[6]) );
  INVX2TS U118 ( .A(n471), .Y(io_byteWrite_8[5]) );
  INVX2TS U119 ( .A(n470), .Y(io_byteWrite_8[4]) );
  INVX2TS U120 ( .A(n469), .Y(io_byteWrite_8[3]) );
  INVX2TS U121 ( .A(n468), .Y(io_byteWrite_8[2]) );
  INVX2TS U122 ( .A(n467), .Y(io_byteWrite_8[1]) );
  INVX2TS U123 ( .A(n466), .Y(io_byteWrite_8[0]) );
  INVX2TS U124 ( .A(n465), .Y(io_byteWrite_9[7]) );
  INVX2TS U125 ( .A(n464), .Y(io_byteWrite_9[6]) );
  INVX2TS U126 ( .A(n463), .Y(io_byteWrite_9[5]) );
  INVX2TS U127 ( .A(n462), .Y(io_byteWrite_9[4]) );
  INVX2TS U128 ( .A(n461), .Y(io_byteWrite_9[3]) );
  INVX2TS U129 ( .A(n460), .Y(io_byteWrite_9[2]) );
  INVX2TS U130 ( .A(n459), .Y(io_byteWrite_9[1]) );
  INVX2TS U131 ( .A(n450), .Y(io_byteWrite_9[0]) );
  INVX2TS U132 ( .A(n457), .Y(io_byteWrite_10[7]) );
  INVX2TS U133 ( .A(n456), .Y(io_byteWrite_10[6]) );
  INVX2TS U134 ( .A(n455), .Y(io_byteWrite_10[5]) );
  INVX2TS U135 ( .A(n454), .Y(io_byteWrite_10[4]) );
  INVX2TS U136 ( .A(n453), .Y(io_byteWrite_10[3]) );
  INVX2TS U137 ( .A(n452), .Y(io_byteWrite_10[2]) );
  INVX2TS U138 ( .A(n451), .Y(io_byteWrite_10[1]) );
  INVX2TS U139 ( .A(n450), .Y(io_byteWrite_10[0]) );
  INVX2TS U140 ( .A(n465), .Y(io_byteWrite_11[7]) );
  INVX2TS U141 ( .A(n464), .Y(io_byteWrite_11[6]) );
  INVX2TS U142 ( .A(n463), .Y(io_byteWrite_11[5]) );
  INVX2TS U143 ( .A(n462), .Y(io_byteWrite_11[4]) );
  INVX2TS U144 ( .A(n461), .Y(io_byteWrite_11[3]) );
  INVX2TS U145 ( .A(n460), .Y(io_byteWrite_11[2]) );
  INVX2TS U146 ( .A(n459), .Y(io_byteWrite_11[1]) );
  INVX2TS U147 ( .A(n458), .Y(io_byteWrite_11[0]) );
  INVX2TS U148 ( .A(n449), .Y(io_byteWrite_12[7]) );
  INVX2TS U149 ( .A(n472), .Y(io_byteWrite_12[6]) );
  INVX2TS U150 ( .A(n471), .Y(io_byteWrite_12[5]) );
  INVX2TS U151 ( .A(n470), .Y(io_byteWrite_12[4]) );
  INVX2TS U152 ( .A(n469), .Y(io_byteWrite_12[3]) );
  INVX2TS U153 ( .A(n468), .Y(io_byteWrite_12[2]) );
  INVX2TS U154 ( .A(n467), .Y(io_byteWrite_12[1]) );
  INVX2TS U155 ( .A(n466), .Y(io_byteWrite_12[0]) );
  INVX2TS U156 ( .A(n449), .Y(io_byteWrite_13[7]) );
  INVX2TS U157 ( .A(n456), .Y(io_byteWrite_13[6]) );
  INVX2TS U158 ( .A(n455), .Y(io_byteWrite_13[5]) );
  INVX2TS U159 ( .A(n454), .Y(io_byteWrite_13[4]) );
  INVX2TS U160 ( .A(n453), .Y(io_byteWrite_13[3]) );
  INVX2TS U161 ( .A(n452), .Y(io_byteWrite_13[2]) );
  INVX2TS U162 ( .A(n451), .Y(io_byteWrite_13[1]) );
  INVX2TS U163 ( .A(n450), .Y(io_byteWrite_13[0]) );
  INVX2TS U164 ( .A(n457), .Y(io_byteWrite_14[7]) );
  INVX2TS U165 ( .A(n456), .Y(io_byteWrite_14[6]) );
  INVX2TS U166 ( .A(n455), .Y(io_byteWrite_14[5]) );
  INVX2TS U167 ( .A(n454), .Y(io_byteWrite_14[4]) );
  INVX2TS U168 ( .A(n453), .Y(io_byteWrite_14[3]) );
  INVX2TS U169 ( .A(n452), .Y(io_byteWrite_14[2]) );
  INVX2TS U170 ( .A(n451), .Y(io_byteWrite_14[1]) );
  INVX2TS U171 ( .A(n458), .Y(io_byteWrite_14[0]) );
  INVX2TS U172 ( .A(n294), .Y(n425) );
  OR2X1TS U173 ( .A(n301), .B(n429), .Y(n278) );
  OR2X1TS U174 ( .A(n301), .B(n426), .Y(n279) );
  NOR2XLTS U175 ( .A(n290), .B(n291), .Y(n280) );
  OR2X1TS U176 ( .A(n445), .B(n435), .Y(n281) );
  OR2X1TS U177 ( .A(n443), .B(n435), .Y(n282) );
  OR2X1TS U178 ( .A(n439), .B(n435), .Y(n283) );
  OR2X1TS U179 ( .A(n445), .B(n429), .Y(n284) );
  OR2X1TS U180 ( .A(n439), .B(n429), .Y(n285) );
  OR2X1TS U181 ( .A(n445), .B(n426), .Y(n286) );
  OR2X1TS U182 ( .A(n443), .B(n426), .Y(n287) );
  OR2X1TS U183 ( .A(n443), .B(n432), .Y(n288) );
  OR2X1TS U184 ( .A(n439), .B(n432), .Y(n289) );
  INVX2TS U185 ( .A(n295), .Y(n298) );
  INVX2TS U186 ( .A(n292), .Y(n297) );
  CLKBUFX2TS U187 ( .A(io_cAddr[2]), .Y(n290) );
  CLKBUFX2TS U188 ( .A(io_cAddr[1]), .Y(n291) );
  INVX2TS U189 ( .A(n280), .Y(n439) );
  CLKBUFX2TS U190 ( .A(io_cAddr[0]), .Y(n292) );
  INVX2TS U191 ( .A(n297), .Y(n302) );
  CLKBUFX2TS U192 ( .A(io_RE), .Y(n293) );
  CLKBUFX2TS U193 ( .A(io_WE), .Y(n294) );
  INVX2TS U194 ( .A(n425), .Y(n438) );
  INVX2TS U195 ( .A(n438), .Y(n304) );
  CLKBUFX2TS U196 ( .A(io_cAddr[3]), .Y(n295) );
  INVX2TS U197 ( .A(n298), .Y(n303) );
  INVX2TS U198 ( .A(n285), .Y(n473) );
  INVX2TS U199 ( .A(n285), .Y(io_bRead[1]) );
  INVX2TS U200 ( .A(n296), .Y(n428) );
  INVX2TS U201 ( .A(n428), .Y(n443) );
  INVX2TS U202 ( .A(n287), .Y(n475) );
  INVX2TS U203 ( .A(n287), .Y(io_bRead[2]) );
  INVX2TS U204 ( .A(n299), .Y(n431) );
  INVX2TS U205 ( .A(n431), .Y(n445) );
  INVX2TS U206 ( .A(n286), .Y(n477) );
  INVX2TS U207 ( .A(n286), .Y(io_bRead[4]) );
  INVX2TS U208 ( .A(n284), .Y(n479) );
  INVX2TS U209 ( .A(n284), .Y(io_bRead[5]) );
  NAND2X1TS U210 ( .A(n290), .B(n291), .Y(n300) );
  INVX2TS U211 ( .A(n300), .Y(n434) );
  INVX2TS U212 ( .A(n434), .Y(n301) );
  INVX2TS U213 ( .A(n279), .Y(n481) );
  INVX2TS U214 ( .A(n279), .Y(io_bRead[6]) );
  INVX2TS U215 ( .A(n278), .Y(n483) );
  INVX2TS U216 ( .A(n278), .Y(io_bRead[7]) );
  INVX2TS U217 ( .A(n283), .Y(n485) );
  INVX2TS U218 ( .A(n283), .Y(io_bRead[8]) );
  INVX2TS U219 ( .A(n289), .Y(n487) );
  INVX2TS U220 ( .A(n289), .Y(io_bRead[9]) );
  INVX2TS U221 ( .A(n282), .Y(n489) );
  INVX2TS U222 ( .A(n282), .Y(io_bRead[10]) );
  INVX2TS U223 ( .A(n288), .Y(n491) );
  INVX2TS U224 ( .A(n288), .Y(io_bRead[11]) );
  INVX2TS U225 ( .A(n281), .Y(n493) );
  INVX2TS U226 ( .A(n281), .Y(io_bRead[12]) );
  CLKBUFX2TS U227 ( .A(io_byteRead_0[7]), .Y(n305) );
  CLKBUFX2TS U228 ( .A(io_byteRead_0[6]), .Y(n306) );
  CLKBUFX2TS U229 ( .A(io_byteRead_0[5]), .Y(n307) );
  CLKBUFX2TS U230 ( .A(io_byteRead_0[4]), .Y(n308) );
  CLKBUFX2TS U231 ( .A(io_byteRead_0[3]), .Y(n309) );
  CLKBUFX2TS U232 ( .A(io_byteRead_0[2]), .Y(n310) );
  CLKBUFX2TS U233 ( .A(io_byteRead_0[1]), .Y(n311) );
  CLKBUFX2TS U234 ( .A(io_byteRead_0[0]), .Y(n312) );
  CLKBUFX2TS U235 ( .A(io_byteRead_1[7]), .Y(n313) );
  CLKBUFX2TS U236 ( .A(io_byteRead_1[6]), .Y(n314) );
  CLKBUFX2TS U237 ( .A(io_byteRead_1[5]), .Y(n315) );
  CLKBUFX2TS U238 ( .A(io_byteRead_1[4]), .Y(n316) );
  CLKBUFX2TS U239 ( .A(io_byteRead_1[3]), .Y(n317) );
  CLKBUFX2TS U240 ( .A(io_byteRead_1[2]), .Y(n318) );
  CLKBUFX2TS U241 ( .A(io_byteRead_1[1]), .Y(n319) );
  CLKBUFX2TS U242 ( .A(io_byteRead_1[0]), .Y(n320) );
  CLKBUFX2TS U243 ( .A(io_byteRead_2[7]), .Y(n321) );
  CLKBUFX2TS U244 ( .A(io_byteRead_2[6]), .Y(n322) );
  CLKBUFX2TS U245 ( .A(io_byteRead_2[5]), .Y(n323) );
  CLKBUFX2TS U246 ( .A(io_byteRead_2[4]), .Y(n324) );
  CLKBUFX2TS U247 ( .A(io_byteRead_2[3]), .Y(n325) );
  CLKBUFX2TS U248 ( .A(io_byteRead_2[2]), .Y(n326) );
  CLKBUFX2TS U249 ( .A(io_byteRead_2[1]), .Y(n327) );
  CLKBUFX2TS U250 ( .A(io_byteRead_2[0]), .Y(n328) );
  CLKBUFX2TS U251 ( .A(io_byteRead_3[7]), .Y(n329) );
  CLKBUFX2TS U252 ( .A(io_byteRead_3[6]), .Y(n330) );
  CLKBUFX2TS U253 ( .A(io_byteRead_3[5]), .Y(n331) );
  CLKBUFX2TS U254 ( .A(io_byteRead_3[4]), .Y(n332) );
  CLKBUFX2TS U255 ( .A(io_byteRead_3[3]), .Y(n333) );
  CLKBUFX2TS U256 ( .A(io_byteRead_3[2]), .Y(n334) );
  CLKBUFX2TS U257 ( .A(io_byteRead_3[1]), .Y(n335) );
  CLKBUFX2TS U258 ( .A(io_byteRead_3[0]), .Y(n336) );
  CLKBUFX2TS U259 ( .A(io_byteRead_4[7]), .Y(n337) );
  CLKBUFX2TS U260 ( .A(io_byteRead_4[6]), .Y(n338) );
  CLKBUFX2TS U261 ( .A(io_byteRead_4[5]), .Y(n339) );
  CLKBUFX2TS U262 ( .A(io_byteRead_4[4]), .Y(n340) );
  CLKBUFX2TS U263 ( .A(io_byteRead_4[3]), .Y(n341) );
  CLKBUFX2TS U264 ( .A(io_byteRead_4[2]), .Y(n342) );
  CLKBUFX2TS U265 ( .A(io_byteRead_4[1]), .Y(n343) );
  CLKBUFX2TS U266 ( .A(io_byteRead_4[0]), .Y(n344) );
  CLKBUFX2TS U267 ( .A(io_byteRead_5[7]), .Y(n345) );
  CLKBUFX2TS U268 ( .A(io_byteRead_5[6]), .Y(n346) );
  CLKBUFX2TS U269 ( .A(io_byteRead_5[5]), .Y(n347) );
  CLKBUFX2TS U270 ( .A(io_byteRead_5[4]), .Y(n348) );
  CLKBUFX2TS U271 ( .A(io_byteRead_5[3]), .Y(n349) );
  CLKBUFX2TS U272 ( .A(io_byteRead_5[2]), .Y(n350) );
  CLKBUFX2TS U273 ( .A(io_byteRead_5[1]), .Y(n351) );
  CLKBUFX2TS U274 ( .A(io_byteRead_5[0]), .Y(n352) );
  CLKBUFX2TS U275 ( .A(io_byteRead_6[7]), .Y(n353) );
  CLKBUFX2TS U276 ( .A(io_byteRead_6[6]), .Y(n354) );
  CLKBUFX2TS U277 ( .A(io_byteRead_6[5]), .Y(n355) );
  CLKBUFX2TS U278 ( .A(io_byteRead_6[4]), .Y(n356) );
  CLKBUFX2TS U279 ( .A(io_byteRead_6[3]), .Y(n357) );
  CLKBUFX2TS U280 ( .A(io_byteRead_6[2]), .Y(n358) );
  CLKBUFX2TS U281 ( .A(io_byteRead_6[1]), .Y(n359) );
  CLKBUFX2TS U282 ( .A(io_byteRead_6[0]), .Y(n360) );
  CLKBUFX2TS U283 ( .A(io_byteRead_7[7]), .Y(n361) );
  CLKBUFX2TS U284 ( .A(io_byteRead_7[6]), .Y(n362) );
  CLKBUFX2TS U285 ( .A(io_byteRead_7[5]), .Y(n363) );
  CLKBUFX2TS U286 ( .A(io_byteRead_7[4]), .Y(n364) );
  CLKBUFX2TS U287 ( .A(io_byteRead_7[3]), .Y(n365) );
  CLKBUFX2TS U288 ( .A(io_byteRead_7[2]), .Y(n366) );
  CLKBUFX2TS U289 ( .A(io_byteRead_7[1]), .Y(n367) );
  CLKBUFX2TS U290 ( .A(io_byteRead_7[0]), .Y(n368) );
  CLKBUFX2TS U291 ( .A(io_byteRead_8[7]), .Y(n369) );
  CLKBUFX2TS U292 ( .A(io_byteRead_8[6]), .Y(n370) );
  CLKBUFX2TS U293 ( .A(io_byteRead_8[5]), .Y(n371) );
  CLKBUFX2TS U294 ( .A(io_byteRead_8[4]), .Y(n372) );
  CLKBUFX2TS U295 ( .A(io_byteRead_8[3]), .Y(n373) );
  CLKBUFX2TS U296 ( .A(io_byteRead_8[2]), .Y(n374) );
  CLKBUFX2TS U297 ( .A(io_byteRead_8[1]), .Y(n375) );
  CLKBUFX2TS U298 ( .A(io_byteRead_8[0]), .Y(n376) );
  CLKBUFX2TS U299 ( .A(io_byteRead_9[7]), .Y(n377) );
  CLKBUFX2TS U300 ( .A(io_byteRead_9[6]), .Y(n378) );
  CLKBUFX2TS U301 ( .A(io_byteRead_9[5]), .Y(n379) );
  CLKBUFX2TS U302 ( .A(io_byteRead_9[4]), .Y(n380) );
  CLKBUFX2TS U303 ( .A(io_byteRead_9[3]), .Y(n381) );
  CLKBUFX2TS U304 ( .A(io_byteRead_9[2]), .Y(n382) );
  CLKBUFX2TS U305 ( .A(io_byteRead_9[1]), .Y(n383) );
  CLKBUFX2TS U306 ( .A(io_byteRead_9[0]), .Y(n384) );
  CLKBUFX2TS U307 ( .A(io_byteRead_10[7]), .Y(n385) );
  CLKBUFX2TS U308 ( .A(io_byteRead_10[6]), .Y(n386) );
  CLKBUFX2TS U309 ( .A(io_byteRead_10[5]), .Y(n387) );
  CLKBUFX2TS U310 ( .A(io_byteRead_10[4]), .Y(n388) );
  CLKBUFX2TS U311 ( .A(io_byteRead_10[3]), .Y(n389) );
  CLKBUFX2TS U312 ( .A(io_byteRead_10[2]), .Y(n390) );
  CLKBUFX2TS U313 ( .A(io_byteRead_10[1]), .Y(n391) );
  CLKBUFX2TS U314 ( .A(io_byteRead_10[0]), .Y(n392) );
  CLKBUFX2TS U315 ( .A(io_byteRead_11[7]), .Y(n393) );
  CLKBUFX2TS U316 ( .A(io_byteRead_11[6]), .Y(n394) );
  CLKBUFX2TS U317 ( .A(io_byteRead_11[5]), .Y(n395) );
  CLKBUFX2TS U318 ( .A(io_byteRead_11[4]), .Y(n396) );
  CLKBUFX2TS U319 ( .A(io_byteRead_11[3]), .Y(n397) );
  CLKBUFX2TS U320 ( .A(io_byteRead_11[2]), .Y(n398) );
  CLKBUFX2TS U321 ( .A(io_byteRead_11[1]), .Y(n399) );
  CLKBUFX2TS U322 ( .A(io_byteRead_11[0]), .Y(n400) );
  CLKBUFX2TS U323 ( .A(io_byteRead_12[7]), .Y(n401) );
  CLKBUFX2TS U324 ( .A(io_byteRead_12[6]), .Y(n402) );
  CLKBUFX2TS U325 ( .A(io_byteRead_12[5]), .Y(n403) );
  CLKBUFX2TS U326 ( .A(io_byteRead_12[4]), .Y(n404) );
  CLKBUFX2TS U327 ( .A(io_byteRead_12[3]), .Y(n405) );
  CLKBUFX2TS U328 ( .A(io_byteRead_12[2]), .Y(n406) );
  CLKBUFX2TS U329 ( .A(io_byteRead_12[1]), .Y(n407) );
  CLKBUFX2TS U330 ( .A(io_byteRead_12[0]), .Y(n408) );
  CLKBUFX2TS U331 ( .A(io_byteRead_13[7]), .Y(n409) );
  CLKBUFX2TS U332 ( .A(io_byteRead_13[6]), .Y(n410) );
  CLKBUFX2TS U333 ( .A(io_byteRead_13[5]), .Y(n411) );
  CLKBUFX2TS U334 ( .A(io_byteRead_13[4]), .Y(n412) );
  CLKBUFX2TS U335 ( .A(io_byteRead_13[3]), .Y(n413) );
  CLKBUFX2TS U336 ( .A(io_byteRead_13[2]), .Y(n414) );
  CLKBUFX2TS U337 ( .A(io_byteRead_13[1]), .Y(n415) );
  CLKBUFX2TS U338 ( .A(io_byteRead_13[0]), .Y(n416) );
  CLKBUFX2TS U339 ( .A(io_byteRead_14[7]), .Y(n417) );
  CLKBUFX2TS U340 ( .A(io_byteRead_14[6]), .Y(n418) );
  CLKBUFX2TS U341 ( .A(io_byteRead_14[5]), .Y(n419) );
  CLKBUFX2TS U342 ( .A(io_byteRead_14[4]), .Y(n420) );
  CLKBUFX2TS U343 ( .A(io_byteRead_14[3]), .Y(n421) );
  CLKBUFX2TS U344 ( .A(io_byteRead_14[2]), .Y(n422) );
  CLKBUFX2TS U345 ( .A(io_byteRead_14[1]), .Y(n423) );
  CLKBUFX2TS U346 ( .A(io_byteRead_14[0]), .Y(n424) );
  INVX2TS U347 ( .A(n425), .Y(n495) );
  INVX2TS U348 ( .A(n425), .Y(n496) );
  INVX2TS U349 ( .A(n280), .Y(n442) );
  OR2X1TS U350 ( .A(n442), .B(n426), .Y(n427) );
  INVX2TS U351 ( .A(n427), .Y(io_bRead[0]) );
  INVX2TS U352 ( .A(n427), .Y(n498) );
  INVX2TS U353 ( .A(n428), .Y(n444) );
  OR2X1TS U354 ( .A(n444), .B(n429), .Y(n430) );
  INVX2TS U355 ( .A(n430), .Y(io_bRead[3]) );
  INVX2TS U356 ( .A(n430), .Y(n500) );
  INVX2TS U357 ( .A(n431), .Y(n447) );
  OR2X1TS U358 ( .A(n447), .B(n432), .Y(n433) );
  INVX2TS U359 ( .A(n433), .Y(io_bRead[13]) );
  INVX2TS U360 ( .A(n433), .Y(n502) );
  OR2X1TS U361 ( .A(n301), .B(n435), .Y(n436) );
  INVX2TS U362 ( .A(n436), .Y(io_bRead[14]) );
  INVX2TS U363 ( .A(n436), .Y(n504) );
  NAND2X1TS U364 ( .A(n438), .B(n437), .Y(n440) );
  NOR2XLTS U365 ( .A(n439), .B(n440), .Y(io_bWrite[0]) );
  NAND3XLTS U366 ( .A(n302), .B(n496), .C(n298), .Y(n441) );
  NOR2XLTS U367 ( .A(n442), .B(n441), .Y(io_bWrite[1]) );
  NOR2XLTS U368 ( .A(n440), .B(n444), .Y(io_bWrite[2]) );
  NOR2XLTS U369 ( .A(n441), .B(n444), .Y(io_bWrite[3]) );
  NOR2XLTS U370 ( .A(n440), .B(n447), .Y(io_bWrite[4]) );
  NOR2XLTS U371 ( .A(n441), .B(n447), .Y(io_bWrite[5]) );
  NOR2XLTS U372 ( .A(n440), .B(n300), .Y(io_bWrite[6]) );
  NOR2XLTS U373 ( .A(n441), .B(n301), .Y(io_bWrite[7]) );
  NAND3XLTS U374 ( .A(n294), .B(n295), .C(n297), .Y(n448) );
  NOR2XLTS U375 ( .A(n442), .B(n448), .Y(io_bWrite[8]) );
  NAND3XLTS U376 ( .A(n495), .B(n292), .C(n303), .Y(n446) );
  NOR2XLTS U377 ( .A(n442), .B(n446), .Y(io_bWrite[9]) );
  NOR2XLTS U378 ( .A(n443), .B(n448), .Y(io_bWrite[10]) );
  NOR2XLTS U379 ( .A(n444), .B(n446), .Y(io_bWrite[11]) );
  NOR2XLTS U380 ( .A(n445), .B(n448), .Y(io_bWrite[12]) );
  NOR2XLTS U381 ( .A(n447), .B(n446), .Y(io_bWrite[13]) );
  NOR2XLTS U382 ( .A(n300), .B(n448), .Y(io_bWrite[14]) );
  INVX2TS U383 ( .A(io_byteWrite_1[7]), .Y(n449) );
  INVX2TS U384 ( .A(io_byteWrite_5[7]), .Y(n457) );
  INVX2TS U385 ( .A(io_byteWrite_1[6]), .Y(n456) );
  INVX2TS U386 ( .A(io_byteWrite_1[5]), .Y(n455) );
  INVX2TS U387 ( .A(io_byteWrite_1[4]), .Y(n454) );
  INVX2TS U388 ( .A(io_byteWrite_1[3]), .Y(n453) );
  INVX2TS U389 ( .A(io_byteWrite_1[2]), .Y(n452) );
  INVX2TS U390 ( .A(io_byteWrite_1[1]), .Y(n451) );
  INVX2TS U391 ( .A(io_byteWrite_1[0]), .Y(n450) );
  INVX2TS U392 ( .A(io_byteWrite_4[7]), .Y(n465) );
  INVX2TS U393 ( .A(io_byteWrite_4[6]), .Y(n464) );
  INVX2TS U394 ( .A(io_byteWrite_4[5]), .Y(n463) );
  INVX2TS U395 ( .A(io_byteWrite_4[4]), .Y(n462) );
  INVX2TS U396 ( .A(io_byteWrite_4[3]), .Y(n461) );
  INVX2TS U397 ( .A(io_byteWrite_4[2]), .Y(n460) );
  INVX2TS U398 ( .A(io_byteWrite_4[1]), .Y(n459) );
  INVX2TS U399 ( .A(io_byteWrite_4[0]), .Y(n458) );
  INVX2TS U400 ( .A(io_byteWrite_3[6]), .Y(n472) );
  INVX2TS U401 ( .A(io_byteWrite_3[5]), .Y(n471) );
  INVX2TS U402 ( .A(io_byteWrite_3[4]), .Y(n470) );
  INVX2TS U403 ( .A(io_byteWrite_3[3]), .Y(n469) );
  INVX2TS U404 ( .A(io_byteWrite_3[2]), .Y(n468) );
  INVX2TS U405 ( .A(io_byteWrite_3[1]), .Y(n467) );
  INVX2TS U406 ( .A(io_byteWrite_3[0]), .Y(n466) );
  INVX2TS U407 ( .A(n505), .Y(io_byteWrite_5[7]) );
  INVX2TS U408 ( .A(n512), .Y(io_byteWrite_4[0]) );
  INVX2TS U409 ( .A(n511), .Y(io_byteWrite_4[1]) );
  INVX2TS U410 ( .A(n510), .Y(io_byteWrite_4[2]) );
  INVX2TS U411 ( .A(n509), .Y(io_byteWrite_4[3]) );
  INVX2TS U412 ( .A(n508), .Y(io_byteWrite_4[4]) );
  INVX2TS U413 ( .A(n507), .Y(io_byteWrite_4[5]) );
  INVX2TS U414 ( .A(n506), .Y(io_byteWrite_4[6]) );
  INVX2TS U415 ( .A(n505), .Y(io_byteWrite_4[7]) );
  INVX2TS U416 ( .A(n512), .Y(io_byteWrite_3[0]) );
  INVX2TS U417 ( .A(n511), .Y(io_byteWrite_3[1]) );
  INVX2TS U418 ( .A(n510), .Y(io_byteWrite_3[2]) );
  INVX2TS U419 ( .A(n509), .Y(io_byteWrite_3[3]) );
  INVX2TS U420 ( .A(n508), .Y(io_byteWrite_3[4]) );
  INVX2TS U421 ( .A(n507), .Y(io_byteWrite_3[5]) );
  INVX2TS U422 ( .A(n506), .Y(io_byteWrite_3[6]) );
  INVX2TS U423 ( .A(n457), .Y(io_byteWrite_3[7]) );
  INVX2TS U424 ( .A(n458), .Y(io_byteWrite_2[0]) );
  INVX2TS U425 ( .A(n459), .Y(io_byteWrite_2[1]) );
  INVX2TS U426 ( .A(n460), .Y(io_byteWrite_2[2]) );
  INVX2TS U427 ( .A(n461), .Y(io_byteWrite_2[3]) );
  INVX2TS U428 ( .A(n462), .Y(io_byteWrite_2[4]) );
  INVX2TS U429 ( .A(n463), .Y(io_byteWrite_2[5]) );
  INVX2TS U430 ( .A(n464), .Y(io_byteWrite_2[6]) );
  INVX2TS U431 ( .A(n465), .Y(io_byteWrite_2[7]) );
  INVX2TS U432 ( .A(n466), .Y(io_byteWrite_0[0]) );
  INVX2TS U433 ( .A(n467), .Y(io_byteWrite_0[1]) );
  INVX2TS U434 ( .A(n468), .Y(io_byteWrite_0[2]) );
  INVX2TS U435 ( .A(n469), .Y(io_byteWrite_0[3]) );
  INVX2TS U436 ( .A(n470), .Y(io_byteWrite_0[4]) );
  INVX2TS U437 ( .A(n471), .Y(io_byteWrite_0[5]) );
  INVX2TS U438 ( .A(n472), .Y(io_byteWrite_0[6]) );
endmodule

